// Copyright (c) 2021 by Rivos Inc.
// Confidential and proprietary, see LICENSE for details.
// SPDX-License-Identifier: LicenseRef-Rivos-Internal-Only


`ifndef DUT_DEFINES

   `define DUT_DEFINES

   `define DUT_READ_SIZE    128
   `define DUT_READ_WORDS   (`DUT_READ_SIZE / 32)
   `define DUT_WRITE_SIZE   288
   `define DUT_WRITE_WORDS  (`DUT_WRITE_SIZE / 32)

`endif
